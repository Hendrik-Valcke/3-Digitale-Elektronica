library IEEE;
use IEEE.std_logic_1164.all;

package LFSRPackage is
  type t_TapsArr is array (integer range <>) of boolean;
end LFSRPackage;
